-- Copyright (C) 2020 Nathan Paul Simons (C2T9uE-code@hardcorehackers.com)
--
-- This program is free software: you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or (at
-- your option) any later version.
--
-- This program is distributed in the hope that it will be useful, but
-- WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
-- General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with this program.  If not, see <http://www.gnu.org/licenses/>.

use std.textio.all;

entity Hello is
end Hello;

architecture Hello_Arch of Hello is

begin  -- Hello_Arch

  p : process
    variable l : line;
  begin
    write(l, String'("Hello, world!"));
    writeline(output, l);
    wait;
  end process;

end Hello_Arch;

-- Local Variables:
--   mode: VHDL
-- End:
-- vi: fileformat=unix expandtab
